module computer



endmodule