module programcounter()

endmodule