`timescale 1ns / 1ns

module testbenchhw5;